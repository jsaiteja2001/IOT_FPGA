----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:53:08 03/11/2024 
-- Design Name: 
-- Module Name:    irmotor - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity irmotor is
Port ( ir : in  STD_LOGIC;
           mot : out  STD_LOGIC);
end irmotor;

architecture Behavioral of irmotor is

begin
process (ir) 
begin 
if ir='0' then 
mot <= '1'; 
else mot <= '0'; 
end if; 
end process; 
end Behavioral;